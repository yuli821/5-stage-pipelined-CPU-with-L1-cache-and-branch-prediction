module BTB_branch_dut_tb();
endmodule : BTB_branch_dut_tb
